module first_program;
   initial
     begin
	$display("Hello Vu");
	$finish;
     end
endmodule
